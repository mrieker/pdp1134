//    Copyright (C) Mike Rieker, Beverly, MA USA
//    www.outerworldapps.com
//
//    This program is free software; you can redistribute it and/or modify
//    it under the terms of the GNU General Public License as published by
//    the Free Software Foundation; version 2 of the License.
//
//    This program is distributed in the hope that it will be useful,
//    but WITHOUT ANY WARRANTY; without even the implied warranty of
//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//    GNU General Public License for more details.
//
//    EXPECT it to FAIL when someone's HeALTh or PROpeRTy is at RISk.
//
//    You should have received a copy of the GNU General Public License
//    along with this program; if not, write to the Free Software
//    Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA
//
//    http://www.gnu.org/licenses/gpl-2.0.html

module synk (input CLOCK, output reg q, input o);
    reg eo, p;
    always @(posedge CLOCK) begin
        if (eo) p <= o;
           else q <= p;
        eo <= ~ eo;
    end
endmodule

// main program for the zynq implementation

module Zynq (
    input  CLOCK,               // 100MHz clock
    input  RESET_N,             // power-on reset

    output LEDoutR,             // IO_B34_LN6 R14
    output LEDoutG,             // IO_B34_LP7 Y16
    output LEDoutB,             // IO_B34_LN7 Y17

    input muxa,                 // multiplexed inputs
    input muxb,
    input muxc,
    input muxd,
    input muxe,
    input muxf,
    input muxh,
    input muxj,
    input muxk,
    input muxl,
    input muxm,
    input muxn,
    input muxp,
    input muxr,
    input muxs,

    output rsel1_h,             // multiplexor selectors
    output rsel2_h,
    output rsel3_h,

    input ac_lo_in_h,           // control inputs
    input bbsy_in_h,
    input dc_lo_in_h,
    input hltgr_in_l,
    input init_in_h,
    input intr_in_h,
    input msyn_in_h,
    input npg_in_l,
    input sack_in_h,
    input ssyn_in_h,

    input[7:4] bg_in_l,         // bus grant inputs

    output reg bbsy_out_h,      // control outputs
    output reg hltrq_out_h,
    output reg init_out_h,
    output reg intr_out_h,
    output reg msyn_out_h,
    output reg npg_out_l,
    output reg npr_out_h,
    output reg pa_out_h,
    output reg pb_out_h,
    output reg sack_out_h,
    output reg ssyn_out_h,

    output reg[17:00] a_out_h,  // address bus outputs
    output reg[7:4]   bg_out_l, // bus grant outputs
    output reg[7:4]   br_out_h, // bus request outputs
    output reg[1:0]   c_out_h,  // control bus outputs
    output reg[15:00] d_out_h,  // data bus outputs

    // arm processor memory bus interface (AXI)
    // we are a slave for accessing the control registers (read and write)
    input[11:00]  saxi_ARADDR,
    output reg    saxi_ARREADY,
    input         saxi_ARVALID,
    input[11:00]  saxi_AWADDR,
    output reg    saxi_AWREADY,
    input         saxi_AWVALID,
    input         saxi_BREADY,
    output[1:0]   saxi_BRESP,
    output reg    saxi_BVALID,
    output[31:00] saxi_RDATA,
    input         saxi_RREADY,
    output[1:0]   saxi_RRESP,
    output reg    saxi_RVALID,
    input[31:00]  saxi_WDATA,
    output reg    saxi_WREADY,
    input         saxi_WVALID);

    // [31:16] = '11'; [15:12] = (log2 len)-1; [11:00] = version
    localparam VERSION = 32'h31314005;

    // bus values that are constants
    assign saxi_BRESP = 0;  // A3.4.4/A10.3 transfer OK
    assign saxi_RRESP = 0;  // A3.4.4/A10.3 transfer OK

    reg[11:02] readaddr, writeaddr;

    reg[55:00] ilaarray[4095:0], ilardata;
    reg[11:00] ilaafter, ilaindex;
    reg ilaarmed;

    ////////////////////////////
    //  internal bus signals  //
    ////////////////////////////

    // _in_ signals: FM_OFF,FM_MAN: zeroes; FM_SIM: from simulator; FM_REAL: from unibus
    // _out_ signals: FM_OFF,FM_MAN: ignored; FM_SIM: to simulator; FM_REAL: to unibus

    reg dev_ac_lo_in_h;
    reg dev_bbsy_in_h;
    reg dev_dc_lo_in_h;
    reg dev_hltgr_in_l;
    reg dev_hltrq_in_h;
    reg dev_intr_in_h;
    reg dev_init_in_h;
    reg dev_msyn_in_h;
    reg dev_msyn_out_h;
    reg dev_npg_in_l;
    reg dev_npg_out_l;
    reg dev_npr_out_h;
    reg dev_sack_in_h;
    reg dev_ssyn_in_h;

    wire dev_hltrq_out_h;
    wire dev_init_out_h;

    reg[1:0] dev_c_in_h;
    reg[1:0] dev_c_out_h;
    reg[7:4] dev_bg_in_l;
    reg[15:00] dev_d_in_h;
    reg[17:00] dev_a_in_h;
    reg[17:00] dev_a_out_h;

    wire dev_bbsy_out_h;
    wire dev_intr_out_h;
    wire dev_sack_out_h;
    wire dev_ssyn_out_h;
    wire[7:4] dev_bg_out_l;
    wire[7:4] dev_br_out_h;
    wire[15:00] dev_d_out_h;

    /////////////////////////////////////////////////////////////
    //  signals coming out of simulator going to internal bus  //
    /////////////////////////////////////////////////////////////

    reg sim_ac_lo_in_h;
    reg sim_bbsy_in_h;
    reg sim_dc_lo_in_h;
    reg sim_hltgr_in_l;
    reg sim_init_in_h;
    reg sim_intr_in_h;
    reg sim_msyn_in_h;
    reg sim_npg_in_l;
    reg sim_sack_in_h;
    reg sim_ssyn_in_h;
    reg[1:0] sim_c_in_h;
    reg[7:4] sim_bg_in_l;
    reg[15:00] sim_d_in_h;
    reg[17:00] sim_a_in_h;

    ///////////////////////////////////////
    //  demultiplex signals from unibus  //
    ///////////////////////////////////////

    // synchronize non-multiplexed signals to fpga clock
    // - worst-case delay of 20nS
    wire syn_ac_lo_in_h, syn_bbsy_in_h, syn_dc_lo_in_h, syn_hltgr_in_l, syn_init_in_h;
    wire syn_intr_in_h, syn_msyn_in_h, syn_npg_in_l, syn_sack_in_h, syn_ssyn_in_h;
    wire[7:4] syn_bg_in_l;
    synk synkac_lo (CLOCK, syn_ac_lo_in_h, ac_lo_in_h);
    synk synkbbsy  (CLOCK, syn_bbsy_in_h,  bbsy_in_h);
    synk synkdc_lo (CLOCK, syn_dc_lo_in_h, dc_lo_in_h);
    synk synkhltgr (CLOCK, syn_hltgr_in_l, hltgr_in_l);
    synk synkinit  (CLOCK, syn_init_in_h,  init_in_h);
    synk synkintr  (CLOCK, syn_intr_in_h,  intr_in_h);
    synk synkmsyn  (CLOCK, syn_msyn_in_h,  msyn_in_h);
    synk synknpg   (CLOCK, syn_npg_in_l,   npg_in_l);
    synk synksack  (CLOCK, syn_sack_in_h,  sack_in_h);
    synk synkssyn  (CLOCK, syn_ssyn_in_h,  ssyn_in_h);
    synk synkbg_4  (CLOCK, syn_bg_in_l[4], bg_in_l[4]);
    synk synkbg_5  (CLOCK, syn_bg_in_l[5], bg_in_l[5]);
    synk synkbg_6  (CLOCK, syn_bg_in_l[6], bg_in_l[6]);
    synk synkbg_7  (CLOCK, syn_bg_in_l[7], bg_in_l[7]);

    // input demux signal latches
    // - loaded from mux pins every 150nS
    reg dmx_hltrq_in_h, dmx_npr_in_h, dmx_pa_in_h, dmx_pb_in_h;
    reg[1:0] dmx_c_in_h;
    reg[7:4] dmx_br_in_h;
    reg[17:00] dmx_a_in_h;
    reg[15:00] dmx_d_in_h;

    // del_msyn_in_h - delayed MUXDELAY*3*10nS so all demuxed signals up-to-date
    // - specifically we care about dmx_a_in_h, dmx_c_in_h, dmx_d_in_h
    //   the other dmx_ signals are just passed to arm for debugging
    localparam MUXDELAY = 15;
    reg del_msyn_in_h;

    reg[5:0] muxcount, muxdelay;
    assign rsel1_h  = muxcount[5:4] == 1;
    assign rsel2_h  = muxcount[5:4] == 2;
    assign rsel3_h  = muxcount[5:4] == 3;

    always @(posedge CLOCK) begin
        if (~ RESET_N) begin
            muxcount <= 8;
        end else begin

            // give transistors 50nS to switch and soak
            if (muxcount[3:0] != MUXDELAY-1) begin
                muxcount[3:0] <= muxcount[3:0] + 1;
            end else begin

                // all soaked in, clock into corresponding flipflops
                if (rsel1_h) begin
                    dmx_pa_in_h    <= muxa;
                    dmx_d_in_h[11] <= muxb;
                    dmx_hltrq_in_h <= muxc;
                    dmx_pb_in_h    <= muxd;
                    dmx_d_in_h[15] <= muxe;
                    dmx_d_in_h[14] <= muxf;
                    dmx_d_in_h[13] <= muxh;
                    dmx_d_in_h[12] <= muxj;
                    dmx_d_in_h[10] <= muxk;
                    dmx_d_in_h[09] <= muxl;
                    dmx_d_in_h[08] <= muxm;
                    dmx_d_in_h[07] <= muxn;
                    dmx_d_in_h[04] <= muxp;
                    dmx_d_in_h[05] <= muxr;
                    dmx_d_in_h[01] <= muxs;
                end
                if (rsel2_h) begin
                    dmx_a_in_h[12] <= muxa;
                    dmx_a_in_h[17] <= muxb;
                    dmx_a_in_h[02] <= muxc;
                    dmx_d_in_h[00] <= muxd;
                    dmx_d_in_h[03] <= muxe;
                    dmx_d_in_h[02] <= muxf;
                    dmx_d_in_h[06] <= muxh;
                    dmx_br_in_h[7] <= muxj;
                    dmx_br_in_h[6] <= muxk;
                    dmx_br_in_h[5] <= muxl;
                    dmx_br_in_h[4] <= muxm;
                    dmx_a_in_h[15] <= muxn;
                    dmx_a_in_h[16] <= muxp;
                    dmx_c_in_h[1]  <= muxr;
                end
                if (rsel3_h) begin
                    dmx_a_in_h[01] <= muxa;
                    dmx_a_in_h[14] <= muxb;
                    dmx_a_in_h[11] <= muxc;
                    dmx_a_in_h[10] <= muxd;
                    dmx_a_in_h[09] <= muxe;
                    dmx_a_in_h[06] <= muxf;
                    dmx_a_in_h[05] <= muxh;
                    dmx_npr_in_h   <= muxj;
                    dmx_a_in_h[00] <= muxk;
                    dmx_c_in_h[0]  <= muxl;
                    dmx_a_in_h[13] <= muxm;
                    dmx_a_in_h[08] <= muxn;
                    dmx_a_in_h[07] <= muxp;
                    dmx_a_in_h[04] <= muxr;
                    dmx_a_in_h[03] <= muxs;
                end

                // increment on to next multiplexor selection
                muxcount[3:0] <= 0;

                // - if FM_MAN mode and non-zero b_rsel_h, use that one
                //   otherwise, cycle on through one to the next
                muxcount[5:4] <=
                    ((regctla[31:30] == FM_MAN) & (regctlb[29:28] != 0)) ? regctlb[29:28] :
                                            (muxcount[5:4] == 3) ? 1 : (muxcount[5:4] + 1);
            end

            // delay msyn_in_h a full demux cycle so we know multiplexed signals are all updated
            // master has given it some delay but give it more to be sure
            if (~ syn_msyn_in_h) begin
                del_msyn_in_h <= 0;                 // drop delayed msyn as soon as external drops
                muxdelay      <= 0;                 // init delay counter for next time
            end else if (muxdelay != MUXDELAY*3-1) begin
                muxdelay      <= muxdelay + 1;
            end else begin                          // see if all 3 clocked in since transition
                del_msyn_in_h <= 1;                 // ok to assert delayed msyn now
            end
        end
    end

    //////////////////////////////////
    //  send signals out to unibus  //
    //////////////////////////////////

    // - hi-Z if OFF or SIM mode
    //   internal bus forwarded to unibus if REAL mode
    //   arm registers forwarded to unibus if MAN mode

    reg[31:00] regctla, regctlb;

    localparam FM_OFF  = 0;
    localparam FM_SIM  = 1;
    localparam FM_REAL = 2;
    localparam FM_MAN  = 3;

    always @(*) begin
        case (regctla[31:30])

            // FM_OFF, FM_SIM
            // - hi-Z all outputs to unibus except forward grant signals on
            // - input muxes shut off
            FM_OFF, FM_SIM: begin
                a_out_h     <= 0;           // sending 0V to gates opens the transistors
                bbsy_out_h  <= 0;
                bg_out_l    <= bg_in_l;     // act as grant jumper card when shut off
                br_out_h    <= 0;
                c_out_h     <= 0;
                d_out_h     <= 0;
                hltrq_out_h <= 0;
                init_out_h  <= 0;
                intr_out_h  <= 0;
                msyn_out_h  <= 0;
                npg_out_l   <= npg_in_l;
                npr_out_h   <= 0;
                pa_out_h    <= 0;
                pb_out_h    <= 0;
                sack_out_h  <= 0;
                ssyn_out_h  <= 0;
            end

            // FM_REAL - forward internal signals out onto unibus
            FM_REAL: begin
                a_out_h     <= dev_a_out_h;
                bbsy_out_h  <= dev_bbsy_out_h;
                bg_out_l    <= dev_bg_out_l;
                br_out_h    <= dev_br_out_h;
                c_out_h     <= dev_c_out_h;
                d_out_h     <= dev_d_out_h;
                hltrq_out_h <= dev_hltrq_out_h;
                init_out_h  <= dev_init_out_h;
                intr_out_h  <= dev_intr_out_h;
                msyn_out_h  <= dev_msyn_out_h;
                npg_out_l   <= dev_npg_out_l;
                npr_out_h   <= dev_npr_out_h;
                pa_out_h    <= 0;
                pb_out_h    <= 0;
                sack_out_h  <= dev_sack_out_h;
                ssyn_out_h  <= dev_ssyn_out_h;
            end

            // FM_MAN - signals come from arm registers
            // - for the grants, =0 passes grant, =1 blocks grant
            FM_MAN: begin
                a_out_h     <= regctlb[17:00];
                bbsy_out_h  <= regctla[26];
                bg_out_l    <= regctlb[27:24] | bg_in_l;
                br_out_h    <= regctlb[23:20];
                c_out_h     <= regctlb[19:18];
                d_out_h     <= regctla[15:00];
                hltrq_out_h <= regctla[25];
                init_out_h  <= regctla[24];
                intr_out_h  <= regctla[23];
                msyn_out_h  <= regctla[22];
                npg_out_l   <= regctla[21]    | npg_in_l;
                npr_out_h   <= regctla[20];
                pa_out_h    <= regctla[19];
                pb_out_h    <= regctla[18];
                sack_out_h  <= regctla[17];
                ssyn_out_h  <= regctla[16];
            end
        endcase
    end

    //////////////////////////////////////////
    //  get input signals for internal bus  //
    //////////////////////////////////////////

    // - zeroes if OFF or MAN
    //   from simulator if SIM
    //   from real unibus if REAL

    always @(*) begin
        case (regctla[31:30])

            // FM_OFF, FM_MAN - zeroes on internal bus
            FM_OFF, FM_MAN: begin
                dev_a_in_h     <= 0;
                dev_ac_lo_in_h <= 0;
                dev_bbsy_in_h  <= 0;
                dev_bg_in_l    <= 15;
                dev_c_in_h     <= 0;
                dev_d_in_h     <= 0;
                dev_dc_lo_in_h <= 0;
                dev_hltgr_in_l <= 1;
                dev_init_in_h  <= ~ RESET_N;
                dev_intr_in_h  <= 0;
                dev_msyn_in_h  <= 0;
                dev_npg_in_l   <= 1;
                dev_sack_in_h  <= 0;
                dev_ssyn_in_h  <= 0;
            end

            // FM_SIM - forward inputs from simulator to internal bus
            FM_SIM: begin
                dev_a_in_h     <= sim_a_in_h;
                dev_ac_lo_in_h <= sim_ac_lo_in_h;
                dev_bbsy_in_h  <= sim_bbsy_in_h;
                dev_bg_in_l    <= sim_bg_in_l;
                dev_c_in_h     <= sim_c_in_h;
                dev_d_in_h     <= sim_d_in_h;
                dev_dc_lo_in_h <= sim_dc_lo_in_h;
                dev_hltgr_in_l <= sim_hltgr_in_l;
                dev_init_in_h  <= sim_init_in_h | ~ RESET_N;
                dev_intr_in_h  <= sim_intr_in_h;
                dev_msyn_in_h  <= sim_msyn_in_h;
                dev_npg_in_l   <= sim_npg_in_l;
                dev_sack_in_h  <= sim_sack_in_h;
                dev_ssyn_in_h  <= sim_ssyn_in_h;
            end

            // FM_REAL - forward inputs from unibus to internal bus
            FM_REAL: begin
                dev_a_in_h     <= dmx_a_in_h;       // demultiplexed
                dev_ac_lo_in_h <= syn_ac_lo_in_h;   // syncd to fpga clock
                dev_bbsy_in_h  <= syn_bbsy_in_h;
                dev_bg_in_l    <= syn_bg_in_l;
                dev_c_in_h     <= dmx_c_in_h;
                dev_d_in_h     <= dmx_d_in_h;
                dev_dc_lo_in_h <= syn_dc_lo_in_h;
                dev_hltgr_in_l <= syn_hltgr_in_l;
                dev_init_in_h  <= syn_init_in_h | ~ RESET_N;
                dev_intr_in_h  <= syn_intr_in_h;
                dev_msyn_in_h  <= del_msyn_in_h;    // delayed until 3 demux cycles complete
                dev_npg_in_l   <= syn_npg_in_l;
                dev_sack_in_h  <= syn_sack_in_h;
                dev_ssyn_in_h  <= syn_ssyn_in_h;
            end
        endcase
    end

    ///////////////////////////////////////////////////////
    //  give arm direct read-only access to unibus pins  //
    ///////////////////////////////////////////////////////

    wire simmode = regctla[31:30] == FM_SIM;

    wire[31:00] regctlc = {
        muxa,               // multiplexed inputs
        muxb,
        muxc,
        muxd,
        muxe,
        muxf,
        muxh,
        muxj,
        muxk,
        muxl,
        muxm,
        muxn,
        muxp,
        muxr,
        muxs,

        rsel1_h,            // multiplexor selectors
        rsel2_h,
        rsel3_h,

        simmode ? sim_ac_lo_in_h : ac_lo_in_h,  // control inputs
        simmode ? sim_bbsy_in_h  : bbsy_in_h,
        simmode ? sim_dc_lo_in_h : dc_lo_in_h,
        simmode ? sim_hltgr_in_l : hltgr_in_l,
        simmode ? sim_init_in_h  : init_in_h,
        simmode ? sim_intr_in_h  : intr_in_h,
        simmode ? sim_msyn_in_h  : msyn_in_h,
        simmode ? sim_npg_in_l   : npg_in_l,
        simmode ? sim_sack_in_h  : sack_in_h,
        simmode ? sim_ssyn_in_h  : ssyn_in_h,

        simmode ? sim_bg_in_l    : bg_in_l      // bus grant inputs
    };

    wire[31:00] regctld = {
        3'b0,

        dev_bbsy_out_h,     // control outputs
        dev_hltrq_out_h,
        dev_init_out_h,
        dev_intr_out_h,
        dev_msyn_out_h,
        dev_npg_out_l,
        dev_npr_out_h,
            pa_out_h,
            pb_out_h,
        dev_sack_out_h,
        dev_ssyn_out_h,

        dev_a_out_h         // address bus outputs
    };

    wire[31:00] regctle = {
        6'b0,

        muxcount,

        simmode ? 1'b0       : dmx_npr_in_h,
        simmode ? 1'b0       : dmx_pa_in_h,
        simmode ? 1'b0       : dmx_pb_in_h,
        simmode ? 1'b0       : dmx_hltrq_in_h,

        simmode ? sim_c_in_h : dmx_c_in_h,
        dev_c_out_h,        // control bus outputs

        simmode ? 1'b0       : dmx_br_in_h,
        dev_br_out_h,       // bus request outputs
        dev_bg_out_l        // bus grant outputs
    };

    wire[31:00] regctlf = {
        14'b0,
        simmode ? sim_a_in_h : dmx_a_in_h
    };

    wire[31:00] regctlg = {
        simmode ? sim_d_in_h : dmx_d_in_h,
        dev_d_out_h         // data bus outputs
    };

    /////////////////////////////////////
    //  arm reading/writing registers  //
    /////////////////////////////////////

    wire[31:00] lmarmrdata, slarmrdata, tt0armrdata;

    assign saxi_RDATA =
        (readaddr        == 10'b0000000000) ? VERSION     :
        (readaddr        == 10'b0000000001) ? regctla     :
        (readaddr        == 10'b0000000010) ? regctlb     :
        (readaddr        == 10'b0000000011) ? regctlc     :
        (readaddr        == 10'b0000000100) ? regctld     :
        (readaddr        == 10'b0000000101) ? regctle     :
        (readaddr        == 10'b0000000110) ? regctlf     :
        (readaddr        == 10'b0000000111) ? regctlg     :
        (readaddr        == 10'b0000010001) ? { ilaarmed, 3'b0, ilaafter, 4'b0, ilaindex } :
        (readaddr        == 10'b0000010010) ? {       ilardata[31:00] } :
        (readaddr        == 10'b0000010011) ? { 8'b0, ilardata[55:32] } :
        (readaddr[11:04] ==  8'b00001000)   ? lmarmrdata  :
        (readaddr[11:04] ==  8'b00001001)   ? slarmrdata  :
        (readaddr[11:04] ==  8'b00001010)   ? tt0armrdata :
        32'hDEADBEEF;

    wire armwrite = saxi_WREADY & saxi_WVALID;              // arm is writing a register (single fpga clock cycle)

    wire lmarmwrite  = armwrite & (writeaddr[11:04] == 8'b00001000);
    wire slarmwrite  = armwrite & (writeaddr[11:04] == 8'b00001001);
    wire tt0armwrite = armwrite & (writeaddr[11:04] == 8'b00001010);

    always @(posedge CLOCK) begin
        if (~ RESET_N) begin
            saxi_ARREADY <= 1;                              // we are ready to accept read address
            saxi_RVALID  <= 0;                              // we are not sending out read data

            saxi_AWREADY <= 1;                              // we are ready to accept write address
            saxi_WREADY  <= 0;                              // we are not ready to accept write data
            saxi_BVALID  <= 0;                              // we are not acknowledging any write

            regctla[31:0] <= FM_OFF;                        // FM_OFF disconnect from bus

        end else begin

            /////////////////////
            //  register read  //
            /////////////////////

            // check for PS sending us a read address
            if (saxi_ARREADY & saxi_ARVALID) begin
                readaddr <= saxi_ARADDR[11:02];             // save address bits we care about
                saxi_ARREADY <= 0;                          // we are no longer accepting a read address
                saxi_RVALID <= 1;                           // we are sending out the corresponding data

            // check for PS acknowledging receipt of data
            end else if (saxi_RVALID & saxi_RREADY) begin
                saxi_ARREADY <= 1;                          // we are ready to accept an address again
                saxi_RVALID <= 0;                           // we are no longer sending out data
            end

            //////////////////////
            //  register write  //
            //////////////////////

            // check for PS sending us write data
            if (armwrite) begin
                case (writeaddr)                            // write data to register
                     10'b0000000001: begin
                        regctla <= saxi_WDATA;
                    end
                    10'b0000000010: begin
                        regctlb <= saxi_WDATA;
                    end
                endcase
                saxi_AWREADY <= 1;                          // we are ready to accept an address again
                saxi_WREADY  <= 0;                          // we are no longer accepting write data
                saxi_BVALID  <= 1;                          // we have accepted the data

            end else begin
                // check for PS sending us a write address
                if (saxi_AWREADY & saxi_AWVALID) begin
                    writeaddr <= saxi_AWADDR[11:02];        // save address bits we care about
                    saxi_AWREADY <= 0;                      // we are no longer accepting a write address
                    saxi_WREADY  <= 1;                      // we are ready to accept write data
                end

                // check for PS acknowledging write acceptance
                if (saxi_BVALID & saxi_BREADY) begin
                    saxi_BVALID <= 0;
                end
            end
        end
    end

    ///////////////
    //  devices  //
    ///////////////

    // little memory
    wire lm_ssyn_out_h;
    wire[15:00] lm_d_out_h;

    lilmem lminst (
        .CLOCK (CLOCK),
        .RESET (~ RESET_N),

        .armraddr (readaddr[3:2]),
        .armrdata (lmarmrdata),
        .armwaddr (writeaddr[3:2]),
        .armwdata (saxi_WDATA),
        .armwrite (lmarmwrite),

        .a_in_h (dev_a_in_h),
        .c_in_h (dev_c_in_h),
        .d_in_h (dev_d_in_h),
        .init_in_h (dev_init_in_h),
        .msyn_in_h (dev_msyn_in_h),

        .d_out_h (lm_d_out_h),
        .ssyn_out_h (lm_ssyn_out_h));

    // switches and lights
    wire sl_sack_out_h, sl_ssyn_out_h;
    wire[15:00] sl_d_out_h;

    swlight slinst (
        .CLOCK (CLOCK),
        .RESET (~ RESET_N),

        .armraddr (readaddr[3:2]),
        .armrdata (slarmrdata),
        .armwaddr (writeaddr[3:2]),
        .armwdata (saxi_WDATA),
        .armwrite (slarmwrite),

        .a_in_h (dev_a_in_h),
        .c_in_h (dev_c_in_h),
        .d_in_h (dev_d_in_h),
        .hltgr_in_l (dev_hltgr_in_l),
        .init_in_h (dev_init_in_h),
        .msyn_in_h (dev_msyn_in_h),

        .d_out_h (sl_d_out_h),
        .hltrq_out_h (dev_hltrq_out_h),
        .init_out_h (dev_init_out_h),
        .sack_out_h (sl_sack_out_h),
        .ssyn_out_h (sl_ssyn_out_h));

    // console tty
    wire tt0intreq, tt0_ssyn_out_h;
    wire[7:0] tt0intvec;
    wire[15:00] tt0_d_out_h;

    dl11 tt0inst (
        .CLOCK (CLOCK),
        .RESET (~ RESET_N),

        .armraddr (readaddr[3:2]),
        .armrdata (tt0armrdata),
        .armwaddr (writeaddr[3:2]),
        .armwdata (saxi_WDATA),
        .armwrite (tt0armwrite),

        .intreq (tt0intreq),
        .intvec (tt0intvec),

        .a_in_h (dev_a_in_h),
        .c_in_h (dev_c_in_h),
        .d_in_h (dev_d_in_h),
        .init_in_h (dev_init_in_h),
        .msyn_in_h (dev_msyn_in_h),

        .d_out_h (tt0_d_out_h),
        .ssyn_out_h (tt0_ssyn_out_h));

    /////////////////////////////
    //  interrupt controllers  //
    /////////////////////////////

    wire[7:0] intvec4 = tt0intreq ? tt0intvec : 1;
    wire[7:0] intvec5 = 1;
    wire[7:0] intvec6 = 1;
    wire[7:0] intvec7 = 1;

    wire irq4_bbsy_out_h, irq4_intr_out_h, irq4_sack_out_h;
    wire irq5_bbsy_out_h, irq5_intr_out_h, irq5_sack_out_h;
    wire irq6_bbsy_out_h, irq6_intr_out_h, irq6_sack_out_h;
    wire irq7_bbsy_out_h, irq7_intr_out_h, irq7_sack_out_h;
    wire[15:00] irq4_d_out_h, irq5_d_out_h, irq6_d_out_h, irq7_d_out_h;

    intctl irq4inst (
        .CLOCK (CLOCK),
        .RESET (dev_init_in_h),

        .intvec (intvec4),

        .bbsy_in_h (dev_bbsy_in_h),
        .bg_in_l   (dev_bg_in_l[4]),
        .sack_in_h (dev_sack_in_h),
        .ssyn_in_h (dev_ssyn_in_h),

        .bbsy_out_h (irq4_bbsy_out_h),
        .bg_out_l   (dev_bg_out_l[4]),
        .br_out_h   (dev_br_out_h[4]),
        .d_out_h    (irq4_d_out_h),
        .intr_out_h (irq4_intr_out_h),
        .sack_out_h (irq4_sack_out_h));

    intctl irq5inst (
        .CLOCK (CLOCK),
        .RESET (dev_init_in_h),

        .intvec (intvec5),

        .bbsy_in_h (dev_bbsy_in_h),
        .bg_in_l   (dev_bg_in_l[5]),
        .sack_in_h (dev_sack_in_h),
        .ssyn_in_h (dev_ssyn_in_h),

        .bbsy_out_h (irq5_bbsy_out_h),
        .bg_out_l   (dev_bg_out_l[5]),
        .br_out_h   (dev_br_out_h[5]),
        .d_out_h    (irq5_d_out_h),
        .intr_out_h (irq5_intr_out_h),
        .sack_out_h (irq5_sack_out_h));

    intctl irq6inst (
        .CLOCK (CLOCK),
        .RESET (dev_init_in_h),

        .intvec (intvec6),

        .bbsy_in_h (dev_bbsy_in_h),
        .bg_in_l   (dev_bg_in_l[6]),
        .sack_in_h (dev_sack_in_h),
        .ssyn_in_h (dev_ssyn_in_h),

        .bbsy_out_h (irq6_bbsy_out_h),
        .bg_out_l   (dev_bg_out_l[6]),
        .br_out_h   (dev_br_out_h[6]),
        .d_out_h    (irq6_d_out_h),
        .intr_out_h (irq6_intr_out_h),
        .sack_out_h (irq6_sack_out_h));

    intctl irq7inst (
        .CLOCK (CLOCK),
        .RESET (dev_init_in_h),

        .intvec (intvec7),

        .bbsy_in_h (dev_bbsy_in_h),
        .bg_in_l   (dev_bg_in_l[7]),
        .sack_in_h (dev_sack_in_h),
        .ssyn_in_h (dev_ssyn_in_h),

        .bbsy_out_h (irq7_bbsy_out_h),
        .bg_out_l   (dev_bg_out_l[7]),
        .br_out_h   (dev_br_out_h[7]),
        .d_out_h    (irq7_d_out_h),
        .intr_out_h (irq7_intr_out_h),
        .sack_out_h (irq7_sack_out_h));

    ////////////////////////////////////////
    //  aggregate all bus output signals  //
    ////////////////////////////////////////

    assign dev_bbsy_out_h = irq4_bbsy_out_h | irq5_bbsy_out_h | irq6_bbsy_out_h | irq7_bbsy_out_h;
    assign dev_d_out_h    = irq4_d_out_h    | irq5_d_out_h    | irq6_d_out_h    | irq7_d_out_h    | lm_d_out_h | sl_d_out_h | tt0_d_out_h;
    assign dev_intr_out_h = irq4_intr_out_h | irq5_intr_out_h | irq6_intr_out_h | irq7_intr_out_h;
    assign dev_sack_out_h = irq4_sack_out_h | irq5_sack_out_h | irq6_sack_out_h | irq7_sack_out_h | sl_sack_out_h;
    assign dev_ssyn_out_h = lm_ssyn_out_h   | sl_ssyn_out_h   | tt0_ssyn_out_h;

    /////////////////////////////////
    //  integrated logic analyzer  //
    /////////////////////////////////

    //  ilaarmed = 0: trigger condition satisfied
    //             1: waiting for trigger condition
    //  ilaafter = number of cycles to record after trigger condition satisfied
    //  ilaindex = next entry in ilaarray to write
    //  iladivid = 0: 100MHz; 1: 50MHz; 2: 33MHz; 4: 25MHz; ...

    reg[3:0] ilacount, iladivid;

    always @(posedge CLOCK) begin
        if (~ RESET_N) begin
            ilaarmed <= 0;
            ilaafter <= 0;
            ilacount <= 0;
            iladivid <= 0;
        end else if (ilacount != iladivid) begin
            ilacount <= ilacount + 1;
        end else begin
            ilacount <= 0;

            if (armwrite & (writeaddr == 10'b0000010001)) begin

                // arm processor is writing control register
                ilaarmed <= saxi_WDATA[31];
                ilaafter <= saxi_WDATA[27:16];
                iladivid <= saxi_WDATA[15:12];
                ilaindex <= saxi_WDATA[11:00];
                ilardata <= ilaarray[saxi_WDATA[11:00]];
            end else begin

                // capture signals while before trigger and for ilaafter cycles thereafter
                if (ilaarmed | (ilaafter != 0)) begin
                    ilaarray[ilaindex] <= {
                        dmx_a_in_h,      // dev_a_in_h,
                            ac_lo_in_h,  // dev_ac_lo_in_h,
                            bbsy_in_h,   // dev_bbsy_in_h,
                            bg_in_l,     // dev_bg_in_l,
                        dmx_br_in_h,     // dev_br_in_h,
                        dmx_c_in_h,      // dev_c_in_h,
                        dmx_d_in_h,      // dev_d_in_h,
                            dc_lo_in_h,  // dev_dc_lo_in_h,
                            hltgr_in_l,  // dev_hltgr_in_l,
                        dmx_hltrq_in_h,  // dev_hltrq_in_h,
                            init_in_h,   // dev_init_in_h,
                            intr_in_h,   // dev_intr_in_h,
                            msyn_in_h,   // dev_msyn_in_h,
                            npg_in_l,    // dev_npg_in_l,
                        dmx_npr_in_h,    // dev_npr_in_h,
                            sack_in_h,   // dev_sack_in_h,
                            ssyn_in_h    // dev_ssyn_in_h
                    };

                    ilaindex <= ilaindex + 1;
                    if (~ ilaarmed) ilaafter <= ilaafter - 1;
                end

                // check trigger condition
                ////if (rsel1_h & muxc) begin   // - hltrq_in_h
                ////if (~ hltgr_in_l) begin
                if (rsel3_h & muxf) begin   // - a_in_h[06]
                    ilaarmed <= 0;
                end
            end
        end
    end
endmodule
