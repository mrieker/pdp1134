//    Copyright (C) Mike Rieker, Beverly, MA USA
//    www.outerworldapps.com
//
//    This program is free software; you can redistribute it and/or modify
//    it under the terms of the GNU General Public License as published by
//    the Free Software Foundation; version 2 of the License.
//
//    This program is distributed in the hope that it will be useful,
//    but WITHOUT ANY WARRANTY; without even the implied warranty of
//    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
//    GNU General Public License for more details.
//
//    EXPECT it to FAIL when someone's HeALTh or PROpeRTy is at RISk.
//
//    You should have received a copy of the GNU General Public License
//    along with this program; if not, write to the Free Software
//    Foundation, Inc., 59 Temple Place, Suite 330, Boston, MA  02111-1307  USA
//
//    http://www.gnu.org/licenses/gpl-2.0.html

// PDP-11 RL01/2 disk interface

module rl11
    #(parameter[17:00] ADDR=18'o774400,
      parameter[7:0] INTVEC=8'o160) (
    input CLOCK, RESET,

    input armwrite,
    input[2:0] armraddr, armwaddr,
    input[31:00] armwdata,
    output[31:00] armrdata,
    output armintrq,

    output reg intreq,
    output[7:0] irvec,
    input intgnt,
    input[7:0] igvec,

    input[17:00] a_in_h,
    input[1:0] c_in_h,
    input[15:00] d_in_h,
    input init_in_h,
    input msyn_in_h,

    output reg[15:00] d_out_h,
    output reg ssyn_out_h

    ,output[15:00] rlcs
    ,output trigger);

    reg enable, fastio, lastready;
    reg[15:00] rlba, rlda, rlmp1, rlmp2, rlmp3;
    reg rlcs_15, rlcs_14, rlcs_00;
    reg[13:01] rlcs_1301;
    reg[3:0] writelocks, writerrors, volchecks, drivetypes, headselects, driveonlines, driveerrors, drivereadys;
    wire[1:0] driveselect = rlcs_1301[09:08];

    assign rlcs = { rlcs_15, rlcs_14, rlcs_1301, rlcs_00 };

    assign armrdata = (armraddr == 0) ? 32'h524C200A : // [31:16] = 'RL'; [15:12] = (log2 nreg) - 1; [11:00] = version
                      (armraddr == 1) ? { rlba,  rlcs  } :
                      (armraddr == 2) ? { rlmp1, rlda  } :
                      (armraddr == 3) ? { rlmp3, rlmp2 } :
                      (armraddr == 4) ? {
                            writelocks,         // 28
                            writerrors,         // 24
                            volchecks,          // 20
                            drivetypes,         // 16
                            headselects,        // 12
                            driveonlines,       // 08
                            driveerrors,        // 04
                            drivereadys } :     // 00
                      (armraddr == 5) ? { enable, fastio, 4'b0, INTVEC, ADDR } :
                      32'hDEADBEEF;

    assign trigger = rlcs_1301[07] & (rlda == 16'o002250);

    assign armintrq = ~ rlcs_1301[07]               // wake z11rl.cc when pdp clears ready bit
                        & (rlcs_1301[03:01] != 0)   //  and neither NOP
                        & (rlcs_1301[03:01] != 2);  //  nor GET STATUS

    assign irvec = INTVEC;

    wire[15:00] rlmpstatus =  {
        2'b0,                       // 15:14
        writelocks[driveselect],    // 13
        2'b0,                       // 12:11
        writerrors[driveselect],    // 10
        volchecks[driveselect],     // 09
        1'b0,                       // 08
        drivetypes[driveselect],    // 07
        headselects[driveselect],   // 06
        1'b0,                       // 05
        driveonlines[driveselect],  // 04
        4'b1101                     // 03:00
    };

    // operate interrupt request
    //  clear either on interrupts disabled or when pdp is reading the vector
    //  set on posedge of ready if interrupts are enabled at the time
    //  - do not interrupt when setting interrupt enable when ready already set
    always @(posedge CLOCK) begin
        if (~ rlcs_1301[07] | ~ rlcs_1301[06] | intgnt & (igvec == irvec)) begin
            intreq <= 0;
        end else if (~ lastready) begin
            intreq <= 1;
        end
        lastready <= rlcs_1301[07];
    end

    // maintain drive ready bit and errors for selected drive
    always @(*) begin
        rlcs_00 = drivereadys[driveselect];
        rlcs_14 = driveerrors[driveselect];
        rlcs_15 = rlcs_14 | rlcs_1301[13] | rlcs_1301[12] | rlcs_1301[11] | rlcs_1301[10];
    end

    // main processing loop
    always @(posedge CLOCK) begin
        if (init_in_h) begin
            if (RESET) begin
                enable <= 0;
                fastio <= 0;
                driveerrors <= 0;
                drivereadys <= 0;
            end

            rlcs_1301   <= 13'b0000001000000;
            rlba[15:00] <= 0;
            rlda[15:00] <= 0;
            d_out_h     <= 0;
            ssyn_out_h  <= 0;
        end

        // arm processor is writing one of the registers
        else if (armwrite) begin
            case (armwaddr)
                1: begin
                    rlba  <= armwdata[31:16];
                    rlcs_1301 <= armwdata[13:01];
                end
                2: begin
                    rlmp1 <= armwdata[31:16];
                    rlda  <= armwdata[15:00];
                end
                3: begin
                    rlmp3 <= armwdata[31:16];
                    rlmp2 <= armwdata[15:00];
                end
                4: begin
                    writelocks   <= armwdata[31:28];
                    writerrors   <= armwdata[27:24];
                    volchecks    <= armwdata[23:20];
                    drivetypes   <= armwdata[19:16];
                    headselects  <= armwdata[15:12];
                    driveonlines <= armwdata[11:08];
                    driveerrors  <= armwdata[07:04];
                    drivereadys  <= armwdata[03:00];
                end
                5: begin
                    enable <= armwdata[31];
                    fastio <= armwdata[30];
                end
            endcase
        end

        // pdp or something else is accessing an i/o register
        else if (~ msyn_in_h & ssyn_out_h) begin
            d_out_h    <= 0;
            ssyn_out_h <= 0;
        end else if (enable & msyn_in_h & (a_in_h[17:03] == ADDR[17:03]) & ~ ssyn_out_h) begin
            ssyn_out_h <= 1;
            if (c_in_h[1]) begin
                case (a_in_h[02:01])

                    // pdp writing control/status register
                    // -    drive select [09:08]
                    //  controller ready [07]     usually cleared so z11rl.cc will process command
                    //  interrupt enable [06]
                    //   bus addr[17:16] [05:04]
                    //     function code [03:01]
                    0: begin
                        if (~ c_in_h[0] |   a_in_h[00]) begin
                            rlcs_1301[09:08] <= d_in_h[09:08];
                        end
                        if (~ c_in_h[0] | ~ a_in_h[00]) begin
                            rlcs_1301[07:01] <= d_in_h[07:01];

                            // see if starting a command
                            if (~ d_in_h[07]) begin

                                // clear error bits if starting any command
                                // this allows rlcs[15] to clear immediately
                                rlcs_1301[13:10] <= 0;

                                // clear drive error bit immediately if GET STATUS with RESET bit
                                // this allows rlcs[15] to clear immediately
                                if ((d_in_h[03:01] == 3'b010) & rlda[03]) begin
                                    driveerrors[d_in_h[09:08]] <= 0;
                                end

                                // clear drive ready immediately when starting a seek
                                if (d_in_h[03:01] == 3'b011) begin
                                    drivereadys[d_in_h[09:08]] <= 0;
                                end
                            end
                        end
                    end

                    // pdp writing bus address
                    1: begin
                        if (~ c_in_h[0] |   a_in_h[00]) begin
                            rlba[15:08] <= d_in_h[15:08];
                        end
                        if (~ c_in_h[0] | ~ a_in_h[00]) begin
                            rlba[07:01] <= d_in_h[07:01];
                        end
                    end

                    // pdp writing disk address
                    2: begin
                        if (~ c_in_h[0] |   a_in_h[00]) begin
                            rlda[15:08] <= d_in_h[15:08];
                        end
                        if (~ c_in_h[0] | ~ a_in_h[00]) begin
                            rlda[07:00] <= d_in_h[07:00];
                        end
                    end

                    // pdp writing multi-purpose
                    3: begin
                        if (~ c_in_h[0] |   a_in_h[00]) begin
                            rlmp1[15:08] <= d_in_h[15:08];
                            rlmp2[15:08] <= d_in_h[15:08];
                            rlmp3[15:08] <= d_in_h[15:08];
                        end
                        if (~ c_in_h[0] | ~ a_in_h[00]) begin
                            rlmp1[07:00] <= d_in_h[07:00];
                            rlmp2[07:00] <= d_in_h[07:00];
                            rlmp3[07:00] <= d_in_h[07:00];
                        end
                    end
                endcase
            end else begin

                // pdp reading a register
                case (a_in_h[02:01])
                    0: begin d_out_h <= rlcs; end
                    1: begin d_out_h <= rlba; end
                    2: begin d_out_h <= rlda; end
                    3: begin d_out_h <= rlmp1; rlmp1 <= rlmp2; rlmp2 <= rlmp3; rlmp3 <= rlmp1; end
                endcase
            end
        end

        // do NOP command here
        else if (~ rlcs_1301[07] & (rlcs_1301[03:01] == 0)) begin
            rlcs_1301[07] <= 1;
        end

        // do GET STATUS command here
        else if (~ rlcs_1301[07] & (rlcs_1301[03:01] == 2)) begin
            if ((rlda[07:00] & 8'o367) != 8'o003) begin
                rlcs_1301[10] <= 1;     // OPI operation incomplete
                rlcs_1301[07] <= 1;
            end else if (rlda[03] & volchecks[driveselect]) begin
                volchecks[driveselect] <= 0;
            end else begin
                rlmp1 <= rlmpstatus;
                rlmp2 <= rlmpstatus;
                rlmp3 <= rlmpstatus;
                rlcs_1301[07] <= 1;
            end
        end
    end
endmodule
